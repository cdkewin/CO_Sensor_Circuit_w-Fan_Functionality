** Profile: "SCHEMATIC1-Performace Analysis"  [ C:\Users\Lenovo\Desktop\final grade cad project\Final Grade CAD Project-PSpiceFiles\SCHEMATIC1\Performace Analysis.sim ] 

** Creating circuit file "Performace Analysis.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\Lenovo\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\23.1.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1000ns 0 
.MC 100 TRAN V([OUT]) YMAX OUTPUT ALL 
.OPTIONS DISTRIBUTION GAUSS
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
