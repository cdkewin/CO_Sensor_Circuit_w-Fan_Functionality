** Profile: "SCHEMATIC1-Monte Carlo"  [ c:\users\lenovo\appdata\roaming\spb_data\cdssetup\workspace\projects\final grade cad project\Final Grade CAD Project-PSpiceFiles\SCHEMATIC1\Monte Carlo.sim ] 

** Creating circuit file "Monte Carlo.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\Lenovo\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\23.1.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1000ns 0 
.MC 10 TRAN V([OUT]) YMAX OUTPUT ALL SEED=200 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
